module AND (
    i1,
    i2,
    out
);

output out;
input i1, i2;

assign out = i1 & i2;

endmodule